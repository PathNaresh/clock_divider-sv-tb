module clk_div(
  input clk,
  input rst,
  output clk_d
);

endmodule
